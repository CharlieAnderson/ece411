module and_gate (

);

endmodule : andgate