import lc3b_types::*;

module decoder (

);

endmodule : decoder 