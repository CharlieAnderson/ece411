module decoder (

);

endmodule : decoder 