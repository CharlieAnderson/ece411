module mp2 (

);


cpu CPU (

);

cache Cache (

);


endmodule : mp2