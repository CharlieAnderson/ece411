module cache (

);



cache_datapath datapath (

);

cache_control controller (

);




endmodule : cache