module or_gate (

);

endmodule : or_gate 